<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="SG Fürth" version="11.69132">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="test" name="Test 6 Bahnen" course="SCM" deadline="2021-05-30" hostclub.url="http://Hier geben Sie Die URL Ihrer Vereinshomepage ein" reservecount="2" result.url="http://Hier die URL für die Live Results Seite" startmethod="1" timing="AUTOMATIC" type="0" state="BY" nation="GER">
      <AGEDATE value="2021-05-30" type="YEAR" />
      <POOL name="Schwimmbad" lanemin="1" lanemax="8" />
      <FACILITY city="test" name="Schwimmbad" nation="GER" state="BY" street="Starsse" zip="12345" />
      <POINTTABLE pointtableid="3011" name="FINA Point Scoring" version="2018" />
      <FEES>
        <FEE type="RELAY" value="1000" />
        <FEE type="LATEENTRY.RELAY" value="500" />
      </FEES>
      <QUALIFY from="2019-06-03" until="1809-06-03" />
      <SESSIONS>
        <SESSION date="2021-06-01" number="1">
          <EVENTS>
            <EVENT eventid="1226" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="1360" number="1" order="1" status="SEEDED" />
                <HEAT heatid="1361" number="2" order="2" status="SEEDED" />
                <HEAT heatid="1362" number="3" order="3" status="SEEDED" />
                <HEAT heatid="1363" number="4" order="4" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1229" gender="F" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="1364" number="1" order="1" status="SEEDED" />
                <HEAT heatid="1365" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1231" gender="M" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <HEATS>
                <HEAT heatid="1366" number="1" order="1" status="SEEDED" />
                <HEAT heatid="1367" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-06-01" number="2">
          <EVENTS>
            <EVENT eventid="1233" gender="F" number="4" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="1368" number="1" order="1" status="SEEDED" />
                <HEAT heatid="1369" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1263" gender="M" number="5" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <HEATS>
                <HEAT heatid="1370" number="1" order="1" status="SEEDED" />
                <HEAT heatid="1371" number="2" order="2" status="SEEDED" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="00003" nation="GER" region="02" clubid="1238" name="SG Tieftaucher">
          <ATHLETES>
            <ATHLETE firstname="Leonie" lastname="Hitzelberger" birthdate="2002-01-01" gender="F" nation="GER" athleteid="1245">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1363" lane="4" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1364" lane="2" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1369" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Siegfried" lastname="Welscher" birthdate="2004-01-01" gender="M" nation="GER" athleteid="1254">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1363" lane="1" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1370" lane="2" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1367" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Dieter" lastname="Zielinski" birthdate="2000-01-01" gender="M" nation="GER" athleteid="1259">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1360" lane="5" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1366" lane="4" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1370" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Gina " lastname="Schimratzki" birthdate="2004-01-01" gender="F" nation="GER" athleteid="1252">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1361" lane="2" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1365" lane="5" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1369" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Joshua " lastname="Wenig" birthdate="2005-01-01" gender="M" nation="GER" athleteid="1239">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1360" lane="3" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1367" lane="1" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1371" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ursula" lastname="Göpel" birthdate="2004-01-01" gender="F" nation="GER" athleteid="1261">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1363" lane="8" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1365" lane="3" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1369" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hendrik" lastname="Lammers" birthdate="2000-01-01" gender="M" nation="GER" athleteid="1247">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1361" lane="4" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1367" lane="6" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1371" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Jochen" lastname="Hartwig" birthdate="2004-01-01" gender="M" nation="GER" athleteid="1251">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1362" lane="8" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1366" lane="2" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1371" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Marlon " lastname="Prigge" birthdate="2003-01-01" gender="F" nation="GER" athleteid="1253">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1363" lane="6" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1364" lane="3" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1369" lane="7" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Torsten" lastname="Roling" birthdate="2003-01-01" gender="M" nation="GER" athleteid="1243">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1362" lane="7" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1367" lane="8" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1370" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Wilma " lastname="Bachmann" birthdate="2004-01-01" gender="F" nation="GER" athleteid="1237">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1360" lane="4" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1365" lane="2" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1368" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Finn" lastname="Rothstein" birthdate="2006-01-01" gender="M" nation="GER" athleteid="1260">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1363" lane="3" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1366" lane="5" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1371" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Lilly " lastname="Hirschochs" birthdate="2005-01-01" gender="F" nation="GER" athleteid="1258">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1362" lane="1" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1365" lane="8" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1368" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Mareike" lastname="Hamann" birthdate="2004-01-01" gender="F" nation="GER" athleteid="1246">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1361" lane="1" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1364" lane="4" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1369" lane="2" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Harry " lastname="Kovacs" birthdate="2001-01-01" gender="M" nation="GER" athleteid="1255">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1361" lane="6" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1367" lane="4" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1370" lane="6" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Ann-Kathrin" lastname="Uzarek" birthdate="2003-01-01" gender="F" nation="GER" athleteid="1244">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1361" lane="3" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1364" lane="6" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1368" lane="6" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00001" nation="GER" region="02" clubid="1236" name="SV Unterwasser">
          <ATHLETES>
            <ATHLETE firstname="Irma" lastname="Herkenhoff" birthdate="2001-01-01" gender="F" nation="GER" athleteid="1240">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1362" lane="3" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1365" lane="7" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1369" lane="8" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Sandra" lastname="Schütte" birthdate="2005-01-01" gender="F" nation="GER" athleteid="1248">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1363" lane="7" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1364" lane="5" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1369" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Hartmut" lastname="Badstuber" birthdate="1998-01-01" gender="M" nation="GER" athleteid="1257">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1361" lane="5" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1366" lane="6" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1371" lane="1" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Tom" lastname="Huppertz" birthdate="1999-01-01" gender="M" nation="GER" athleteid="1256">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1363" lane="2" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1371" lane="4" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1367" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Evelyn" lastname="Gustenberg" birthdate="2005-01-01" gender="F" nation="GER" athleteid="1250">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1363" lane="5" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1365" lane="4" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1368" lane="4" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Matthias " lastname="Rumpel" birthdate="2004-01-01" gender="M" nation="GER" athleteid="1249">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1361" lane="7" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1366" lane="3" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1370" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Rita " lastname="Fröse" birthdate="2008-01-01" gender="F" nation="GER" athleteid="1235">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1362" lane="4" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1365" lane="6" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1368" lane="3" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Steffen" lastname="Olbertz" birthdate="2004-01-01" gender="M" nation="GER" athleteid="1241">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1362" lane="2" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1367" lane="7" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1371" lane="7" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Erna " lastname="Birk" birthdate="2002-01-01" gender="F" nation="GER" athleteid="1242">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1362" lane="5" />
                <ENTRY entrytime="NT" eventid="1229" heatid="1365" lane="1" />
                <ENTRY entrytime="NT" eventid="1233" heatid="1369" lane="5" />
              </ENTRIES>
            </ATHLETE>
            <ATHLETE firstname="Günther" lastname="Hartz" birthdate="1996-01-01" gender="M" nation="GER" athleteid="1262">
              <ENTRIES>
                <ENTRY entrytime="NT" eventid="1226" heatid="1362" lane="6" />
                <ENTRY entrytime="NT" eventid="1231" heatid="1367" lane="2" />
                <ENTRY entrytime="NT" eventid="1263" heatid="1371" lane="5" />
              </ENTRIES>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
